module InstructionMemory
#(parameter Inst_Num = 150, parameter Inst_Num_BIT = 8)
(Inst_Address, Instruction);
	input [Inst_Num_BIT - 1:0] Inst_Address;
	output reg [31:0] Instruction;

	always @ (*)begin
		case(Inst_Address)
			'd0:	Instruction <= 32'b00111100000000010110000101100101;
			'd1:	Instruction <= 32'b00110100001000010110000101100101;
			'd2:	Instruction <= 32'b00000000000000010100000000100000;
			'd3:	Instruction <= 32'b10101100000010000000000000000000;
			'd4:	Instruction <= 32'b10101100000010000000000000000100;
			'd5:	Instruction <= 32'b00100000000010000110000101100101;
			'd6:	Instruction <= 32'b10101100000010000000000000001000;
			'd7:	Instruction <= 32'b00100000000010000110010101100001;
			'd8:	Instruction <= 32'b10101100000010000000001000000000;
			'd9:	Instruction <= 32'b00100000000001000000000000001010;
			'd10:	Instruction <= 32'b00100000000001010000000000000000;
			'd11:	Instruction <= 32'b00100000000001100000000000000010;
			'd12:	Instruction <= 32'b00100000000001110000001000000000;
			'd13:	Instruction <= 32'b00001100000000000000000001110111;
			'd14:	Instruction <= 32'b00100000000010000000000000000001;
			'd15:	Instruction <= 32'b00111100000000010100000000000000;
			'd16:	Instruction <= 32'b00000000001000000000100000100001;
			'd17:	Instruction <= 32'b10101100001010000000000000001100;
			'd18:	Instruction <= 32'b00111100000000010000000011111111;
			'd19:	Instruction <= 32'b00110100001000011111111111111111;
			'd20:	Instruction <= 32'b00000000000000010100000000100001;
			'd21:	Instruction <= 32'b00010001000000000000000000000010;
			'd22:	Instruction <= 32'b00100001000010001111111111111111;
			'd23:	Instruction <= 32'b00001000000000000000000000010101;
			'd24:	Instruction <= 32'b00100000000010000000000000000011;
			'd25:	Instruction <= 32'b00111100000000010100000000000000;
			'd26:	Instruction <= 32'b00000000001000000000100000100001;
			'd27:	Instruction <= 32'b10101100001010000000000000001100;
			'd28:	Instruction <= 32'b00000000000000100010000000100001;
			'd29:	Instruction <= 32'b00111100000000010100000000000000;
			'd30:	Instruction <= 32'b00110100001000010000000000010000;
			'd31:	Instruction <= 32'b00000000000000011000000000100000;
			'd32:	Instruction <= 32'b00000000000000101000100000100001;
			'd33:	Instruction <= 32'b00100000000100100000000000010000;
			'd34:	Instruction <= 32'b00000000000100101001000001000010;
			'd35:	Instruction <= 32'b00010110010000000000000000000001;
			'd36:	Instruction <= 32'b00100000000100100000000000001000;
			'd37:	Instruction <= 32'b00100100000010000010011100010000;
			'd38:	Instruction <= 32'b00010001000000000000000000000010;
			'd39:	Instruction <= 32'b00100001000010001111111111111111;
			'd40:	Instruction <= 32'b00001000000000000000000000100110;
			'd41:	Instruction <= 32'b00000000000100100001001000000000;
			'd42:	Instruction <= 32'b00100000000000010000000000000001;
			'd43:	Instruction <= 32'b00010000001100100000000000001010;
			'd44:	Instruction <= 32'b00100000000000010000000000000010;
			'd45:	Instruction <= 32'b00010000001100100000000000000110;
			'd46:	Instruction <= 32'b00100000000000010000000000000100;
			'd47:	Instruction <= 32'b00010000001100100000000000000010;
			'd48:	Instruction <= 32'b00000000000001000100010000000000;
			'd49:	Instruction <= 32'b00001000000000000000000000110111;
			'd50:	Instruction <= 32'b00000000000001000100010100000000;
			'd51:	Instruction <= 32'b00001000000000000000000000110111;
			'd52:	Instruction <= 32'b00000000000001000100011000000000;
			'd53:	Instruction <= 32'b00001000000000000000000000110111;
			'd54:	Instruction <= 32'b00000000000001000100011100000000;
			'd55:	Instruction <= 32'b00000000000010000100011100000010;
			'd56:	Instruction <= 32'b00100000000000010000000000000000;
			'd57:	Instruction <= 32'b00010000001010000000000000111010;
			'd58:	Instruction <= 32'b00100000000000010000000000000001;
			'd59:	Instruction <= 32'b00010000001010000000000000110110;
			'd60:	Instruction <= 32'b00100000000000010000000000000010;
			'd61:	Instruction <= 32'b00010000001010000000000000110010;
			'd62:	Instruction <= 32'b00100000000000010000000000000011;
			'd63:	Instruction <= 32'b00010000001010000000000000101110;
			'd64:	Instruction <= 32'b00100000000000010000000000000100;
			'd65:	Instruction <= 32'b00010000001010000000000000101010;
			'd66:	Instruction <= 32'b00100000000000010000000000000101;
			'd67:	Instruction <= 32'b00010000001010000000000000100110;
			'd68:	Instruction <= 32'b00100000000000010000000000000110;
			'd69:	Instruction <= 32'b00010000001010000000000000100010;
			'd70:	Instruction <= 32'b00100000000000010000000000000111;
			'd71:	Instruction <= 32'b00010000001010000000000000011110;
			'd72:	Instruction <= 32'b00100000000000010000000000001000;
			'd73:	Instruction <= 32'b00010000001010000000000000011010;
			'd74:	Instruction <= 32'b00100000000000010000000000001001;
			'd75:	Instruction <= 32'b00010000001010000000000000010110;
			'd76:	Instruction <= 32'b00100000000000010000000000001010;
			'd77:	Instruction <= 32'b00010000001010000000000000010010;
			'd78:	Instruction <= 32'b00100000000000010000000000001011;
			'd79:	Instruction <= 32'b00010000001010000000000000001110;
			'd80:	Instruction <= 32'b00100000000000010000000000001100;
			'd81:	Instruction <= 32'b00010000001010000000000000001010;
			'd82:	Instruction <= 32'b00100000000000010000000000001101;
			'd83:	Instruction <= 32'b00010000001010000000000000000110;
			'd84:	Instruction <= 32'b00100000000000010000000000001110;
			'd85:	Instruction <= 32'b00010000001010000000000000000010;
			'd86:	Instruction <= 32'b00100000010000100000000001110001;
			'd87:	Instruction <= 32'b00001000000000000000000001110101;
			'd88:	Instruction <= 32'b00100000010000100000000001111001;
			'd89:	Instruction <= 32'b00001000000000000000000001110101;
			'd90:	Instruction <= 32'b00100000010000100000000001011110;
			'd91:	Instruction <= 32'b00001000000000000000000001110101;
			'd92:	Instruction <= 32'b00100000010000100000000000111001;
			'd93:	Instruction <= 32'b00001000000000000000000001110101;
			'd94:	Instruction <= 32'b00100000010000100000000001111100;
			'd95:	Instruction <= 32'b00001000000000000000000001110101;
			'd96:	Instruction <= 32'b00100000010000100000000001110111;
			'd97:	Instruction <= 32'b00001000000000000000000001110101;
			'd98:	Instruction <= 32'b00100000010000100000000001101111;
			'd99:	Instruction <= 32'b00001000000000000000000001110101;
			'd100:	Instruction <= 32'b00100000010000100000000001111111;
			'd101:	Instruction <= 32'b00001000000000000000000001110101;
			'd102:	Instruction <= 32'b00100000010000100000000000000111;
			'd103:	Instruction <= 32'b00001000000000000000000001110101;
			'd104:	Instruction <= 32'b00100000010000100000000001111101;
			'd105:	Instruction <= 32'b00001000000000000000000001110101;
			'd106:	Instruction <= 32'b00100000010000100000000001101101;
			'd107:	Instruction <= 32'b00001000000000000000000001110101;
			'd108:	Instruction <= 32'b00100000010000100000000001100110;
			'd109:	Instruction <= 32'b00001000000000000000000001110101;
			'd110:	Instruction <= 32'b00100000010000100000000001001111;
			'd111:	Instruction <= 32'b00001000000000000000000001110101;
			'd112:	Instruction <= 32'b00100000010000100000000001011011;
			'd113:	Instruction <= 32'b00001000000000000000000001110101;
			'd114:	Instruction <= 32'b00100000010000100000000000000110;
			'd115:	Instruction <= 32'b00001000000000000000000001110101;
			'd116:	Instruction <= 32'b00100000010000100000000000111111;
			'd117:	Instruction <= 32'b10101110000000100000000000000000;
			'd118:	Instruction <= 32'b00001000000000000000000000100010;
			'd119:	Instruction <= 32'b00100011101111011111111111110100;
			'd120:	Instruction <= 32'b10101111101111110000000000001000;
			'd121:	Instruction <= 32'b10101111101100000000000000000100;
			'd122:	Instruction <= 32'b10101111101100010000000000000000;
			'd123:	Instruction <= 32'b00000000100001101000000000100010;
			'd124:	Instruction <= 32'b00000000000001101000100000100001;
			'd125:	Instruction <= 32'b00100100000010100000000000000000;
			'd126:	Instruction <= 32'b00100100000010000000000000000000;
			'd127:	Instruction <= 32'b00000010000010000000100000101010;
			'd128:	Instruction <= 32'b00010100001000000000000000001111;
			'd129:	Instruction <= 32'b00100100000010010000000000000000;
			'd130:	Instruction <= 32'b00000001001100010000100000101010;
			'd131:	Instruction <= 32'b00010000001000000000000000001000;
			'd132:	Instruction <= 32'b00000001000010010101100000100000;
			'd133:	Instruction <= 32'b00000000101010110101100000100000;
			'd134:	Instruction <= 32'b10010001011010110000000000000000;
			'd135:	Instruction <= 32'b00000000111010010110000000100000;
			'd136:	Instruction <= 32'b10010001100011000000000000000000;
			'd137:	Instruction <= 32'b00010101011011000000000000000010;
			'd138:	Instruction <= 32'b00100001001010010000000000000001;
			'd139:	Instruction <= 32'b00001000000000000000000010000010;
			'd140:	Instruction <= 32'b00010101001100010000000000000001;
			'd141:	Instruction <= 32'b00100001010010100000000000000001;
			'd142:	Instruction <= 32'b00100001000010000000000000000001;
			'd143:	Instruction <= 32'b00001000000000000000000001111111;
			'd144:	Instruction <= 32'b00000000000010100001000000100001;
			'd145:	Instruction <= 32'b10001111101111110000000000001000;
			'd146:	Instruction <= 32'b10001111101100000000000000000100;
			'd147:	Instruction <= 32'b10001111101100010000000000000000;
			'd148:	Instruction <= 32'b00100011101111010000000000001100;
			'd149:	Instruction <= 32'b00000011111000000000000000001000;
			default: Instruction <= 32'h00000000;
		endcase
	end
endmodule
module InstructionMemory
#(parameter Inst_Num = 46, parameter Inst_Num_BIT = 8)
(Inst_Address, Instruction);
	input [Inst_Num_BIT-1:0] Inst_Address;
	output reg [31:0] Instruction;

	always @ (*)begin
		case(Inst_Address)
			'd0:	Instruction <= 32'b00111100000000010110000101100101;
			'd1:	Instruction <= 32'b00110100001000010110000101100101;
			'd2:	Instruction <= 32'b00000000000000010100000000100000;
			'd3:	Instruction <= 32'b10101100000010000000000000000000;
			'd4:	Instruction <= 32'b10101100000010000000000000000100;
			'd5:	Instruction <= 32'b00100000000010000110000101100101;
			'd6:	Instruction <= 32'b10101100000010000000000000001000;
			'd7:	Instruction <= 32'b00100000000010000110010101100001;
			'd8:	Instruction <= 32'b10101100000010000000001000000000;
			'd9:	Instruction <= 32'b00100000000001000000000000001010;
			'd10:	Instruction <= 32'b00100000000001010000000000000000;
			'd11:	Instruction <= 32'b00100000000001100000000000000010;
			'd12:	Instruction <= 32'b00100000000001110000001000000000;
			'd13:	Instruction <= 32'b00001100000000000000000000001111;
			'd14:	Instruction <= 32'b00001000000000000000000000001110;
			'd15:	Instruction <= 32'b00100011101111011111111111110100;
			'd16:	Instruction <= 32'b10101111101111110000000000001000;
			'd17:	Instruction <= 32'b10101111101100000000000000000100;
			'd18:	Instruction <= 32'b10101111101100010000000000000000;
			'd19:	Instruction <= 32'b00000000100001101000000000100010;
			'd20:	Instruction <= 32'b00000000000001101000100000100001;
			'd21:	Instruction <= 32'b00100100000010100000000000000000;
			'd22:	Instruction <= 32'b00100100000010000000000000000000;
			'd23:	Instruction <= 32'b00000010000010000000100000101010;
			'd24:	Instruction <= 32'b00010100001000000000000000001111;
			'd25:	Instruction <= 32'b00100100000010010000000000000000;
			'd26:	Instruction <= 32'b00000001001100010000100000101010;
			'd27:	Instruction <= 32'b00010000001000000000000000001000;
			'd28:	Instruction <= 32'b00000001000010010101100000100000;
			'd29:	Instruction <= 32'b00000000101010110101100000100000;
			'd30:	Instruction <= 32'b10010001011010110000000000000000;
			'd31:	Instruction <= 32'b00000000111010010110000000100000;
			'd32:	Instruction <= 32'b10010001100011000000000000000000;
			'd33:	Instruction <= 32'b00010101011011000000000000000010;
			'd34:	Instruction <= 32'b00100001001010010000000000000001;
			'd35:	Instruction <= 32'b00001000000000000000000000011010;
			'd36:	Instruction <= 32'b00010101001100010000000000000001;
			'd37:	Instruction <= 32'b00100001010010100000000000000001;
			'd38:	Instruction <= 32'b00100001000010000000000000000001;
			'd39:	Instruction <= 32'b00001000000000000000000000010111;
			'd40:	Instruction <= 32'b00000000000010100001000000100001;
			'd41:	Instruction <= 32'b10001111101111110000000000001000;
			'd42:	Instruction <= 32'b10001111101100000000000000000100;
			'd43:	Instruction <= 32'b10001111101100010000000000000000;
			'd44:	Instruction <= 32'b00100011101111010000000000001100;
			'd45:	Instruction <= 32'b00000011111000000000000000001000;
			default: Instruction <= 32'h00000000;
		endcase
	end
endmodule